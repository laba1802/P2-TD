`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:10:43 03/21/2017 
// Design Name: 
// Module Name:    comparatorQueue 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module comparatorQueue(
    input [2:0] floorCall,
    input [2:0] actualState,
    input [2:0] firstPosMem,
    input up_down_actual,
    input up_down_call
    );

	//always @ (floorCall)

endmodule
